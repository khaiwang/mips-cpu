`timescale 1ns / 1ns
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/10/15 20:28:59
// Design Name: 
// Module Name: alu
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module Adder_32(input [31:0] A, input [31:0] B, input cin, output [31:0] sum, output Over);
    wire [31:0] c, p, g;
    assign p = A ^ B;
    assign g = A & B;
    assign c[0] = g[0]| (cin & p[0]);
    assign c[1] = g[1] | (p[1] & g[0])| (cin & p[0] & p[1]);
    assign c[2] = g[2] | (p[2] & g[1]) | (p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2]);
    assign c[3] = g[3] | (p[3] & g[2]) | (p[3] & p[2] & g[1]) | (p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3]);
    assign c[4] = g[4] | (p[4] & g[3]) | (p[4] & p[3] & g[2]) | (p[4] & p[3] & p[2] & g[1]) | (p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4]);
    assign c[5] = g[5] | (p[5] & g[4]) | (p[5] & p[4] & g[3]) | (p[5] & p[4] & p[3] & g[2]) | (p[5] & p[4] & p[3] & p[2] & g[1]) | (p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5]);
    assign c[6] = g[6] | (p[6] & g[5]) | (p[6] & p[5] & g[4]) | (p[6] & p[5] & p[4] & g[3]) | (p[6] & p[5] & p[4] & p[3] & g[2]) | (p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6]);
    assign c[7] = g[7] | (p[7] & g[6]) | (p[7] & p[6] & g[5]) | (p[7] & p[6] & p[5] & g[4]) | (p[7] & p[6] & p[5] & p[4] & g[3]) | (p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7]);
    assign c[8] = g[8] | (p[8] & g[7]) | (p[8] & p[7] & g[6]) | (p[8] & p[7] & p[6] & g[5]) | (p[8] & p[7] & p[6] & p[5] & g[4]) | (p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8]);
    assign c[9] = g[9] | (p[9] & g[8]) | (p[9] & p[8] & g[7]) | (p[9] & p[8] & p[7] & g[6]) | (p[9] & p[8] & p[7] & p[6] & g[5]) | (p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9]);
    assign c[10] = g[10] | (p[10] & g[9]) | (p[10] & p[9] & g[8]) | (p[10] & p[9] & p[8] & g[7]) | (p[10] & p[9] & p[8] & p[7] & g[6]) | (p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10]);
    assign c[11] = g[11] | (p[11] & g[10]) | (p[11] & p[10] & g[9]) | (p[11] & p[10] & p[9] & g[8]) | (p[11] & p[10] & p[9] & p[8] & g[7]) | (p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11]);
    assign c[12] = g[12] | (p[12] & g[11]) | (p[12] & p[11] & g[10]) | (p[12] & p[11] & p[10] & g[9]) | (p[12] & p[11] & p[10] & p[9] & g[8]) | (p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12]);
    assign c[13] = g[13] | (p[13] & g[12]) | (p[13] & p[12] & g[11]) | (p[13] & p[12] & p[11] & g[10]) | (p[13] & p[12] & p[11] & p[10] & g[9]) | (p[13] & p[12] & p[11] & p[10] & p[9] & g[8]) | (p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13]);
    assign c[14] = g[14] | (p[14] & g[13]) | (p[14] & p[13] & g[12]) | (p[14] & p[13] & p[12] & g[11]) | (p[14] & p[13] & p[12] & p[11] & g[10]) | (p[14] & p[13] & p[12] & p[11] & p[10] & g[9]) | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8]) | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14]);
    assign c[15] = g[15] | (p[15] & g[14]) | (p[15] & p[14] & g[13]) | (p[15] & p[14] & p[13] & g[12]) | (p[15] & p[14] & p[13] & p[12] & g[11]) | (p[15] & p[14] & p[13] & p[12] & p[11] & g[10]) | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9]) | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8]) | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15]);
    assign c[16] = g[16] | (p[16] & g[15]) | (p[16] & p[15] & g[14]) | (p[16] & p[15] & p[14] & g[13]) | (p[16] & p[15] & p[14] & p[13] & g[12]) | (p[16] & p[15] & p[14] & p[13] & p[12] & g[11]) | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10]) | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9]) | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8]) | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16]);
    assign c[17] = g[17] | (p[17] & g[16]) | (p[17] & p[16] & g[15]) | (p[17] & p[16] & p[15] & g[14]) | (p[17] & p[16] & p[15] & p[14] & g[13]) | (p[17] & p[16] & p[15] & p[14] & p[13] & g[12]) | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11]) | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10]) | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9]) | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8]) | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17]);
    assign c[18] = g[18] | (p[18] & g[17]) | (p[18] & p[17] & g[16]) | (p[18] & p[17] & p[16] & g[15]) | (p[18] & p[17] & p[16] & p[15] & g[14]) | (p[18] & p[17] & p[16] & p[15] & p[14] & g[13]) | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12]) | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11]) | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10]) | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9]) | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8]) | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18]);
    assign c[19] = g[19] | (p[19] & g[18]) | (p[19] & p[18] & g[17]) | (p[19] & p[18] & p[17] & g[16]) | (p[19] & p[18] & p[17] & p[16] & g[15]) | (p[19] & p[18] & p[17] & p[16] & p[15] & g[14]) | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13]) | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12]) | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11]) | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10]) | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9]) | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8]) | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19]);
    assign c[20] = g[20] | (p[20] & g[19]) | (p[20] & p[19] & g[18]) | (p[20] & p[19] & p[18] & g[17]) | (p[20] & p[19] & p[18] & p[17] & g[16]) | (p[20] & p[19] & p[18] & p[17] & p[16] & g[15]) | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14]) | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13]) | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12]) | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11]) | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10]) | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9]) | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8]) | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20]);
    assign c[21] = g[21] | (p[21] & g[20]) | (p[21] & p[20] & g[19]) | (p[21] & p[20] & p[19] & g[18]) | (p[21] & p[20] & p[19] & p[18] & g[17]) | (p[21] & p[20] & p[19] & p[18] & p[17] & g[16]) | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15]) | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14]) | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13]) | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12]) | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11]) | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10]) | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9]) | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8]) | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21]);
    assign c[22] = g[22] | (p[22] & g[21]) | (p[22] & p[21] & g[20]) | (p[22] & p[21] & p[20] & g[19]) | (p[22] & p[21] & p[20] & p[19] & g[18]) | (p[22] & p[21] & p[20] & p[19] & p[18] & g[17]) | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & g[16]) | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15]) | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14]) | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13]) | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12]) | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11]) | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10]) | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9]) | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8]) | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22]);
    assign c[23] = g[23] | (p[23] & g[22]) | (p[23] & p[22] & g[21]) | (p[23] & p[22] & p[21] & g[20]) | (p[23] & p[22] & p[21] & p[20] & g[19]) | (p[23] & p[22] & p[21] & p[20] & p[19] & g[18]) | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & g[17]) | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & g[16]) | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15]) | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14]) | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13]) | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12]) | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11]) | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10]) | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9]) | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8]) | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23]);
    assign c[24] = g[24] | (p[24] & g[23]) | (p[24] & p[23] & g[22]) | (p[24] & p[23] & p[22] & g[21]) | (p[24] & p[23] & p[22] & p[21] & g[20]) | (p[24] & p[23] & p[22] & p[21] & p[20] & g[19]) | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & g[18]) | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & g[17]) | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & g[16]) | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15]) | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14]) | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13]) | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12]) | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11]) | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10]) | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9]) | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8]) | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24]);
    assign c[25] = g[25] | (p[25] & g[24]) | (p[25] & p[24] & g[23]) | (p[25] & p[24] & p[23] & g[22]) | (p[25] & p[24] & p[23] & p[22] & g[21]) | (p[25] & p[24] & p[23] & p[22] & p[21] & g[20]) | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & g[19]) | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & g[18]) | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & g[17]) | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & g[16]) | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15]) | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14]) | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13]) | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12]) | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11]) | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10]) | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9]) | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8]) | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25]);
    assign c[26] = g[26] | (p[26] & g[25]) | (p[26] & p[25] & g[24]) | (p[26] & p[25] & p[24] & g[23]) | (p[26] & p[25] & p[24] & p[23] & g[22]) | (p[26] & p[25] & p[24] & p[23] & p[22] & g[21]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & g[20]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & g[19]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & g[18]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & g[17]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & g[16]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26]);
    assign c[27] = g[27] | (p[27] & g[26]) | (p[27] & p[26] & g[25]) | (p[27] & p[26] & p[25] & g[24]) | (p[27] & p[26] & p[25] & p[24] & g[23]) | (p[27] & p[26] & p[25] & p[24] & p[23] & g[22]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & g[21]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & g[20]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & g[19]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & g[18]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & g[17]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & g[16]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27]);
    assign c[28] = g[28] | (p[28] & g[27]) | (p[28] & p[27] & g[26]) | (p[28] & p[27] & p[26] & g[25]) | (p[28] & p[27] & p[26] & p[25] & g[24]) | (p[28] & p[27] & p[26] & p[25] & p[24] & g[23]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & g[22]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & g[21]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & g[20]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & g[19]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & g[18]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & g[17]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & g[16]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28]);
    assign c[29] = g[29] | (p[29] & g[28]) | (p[29] & p[28] & g[27]) | (p[29] & p[28] & p[27] & g[26]) | (p[29] & p[28] & p[27] & p[26] & g[25]) | (p[29] & p[28] & p[27] & p[26] & p[25] & g[24]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & g[23]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & g[22]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & g[21]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & g[20]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & g[19]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & g[18]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & g[17]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & g[16]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29]);
    assign c[30] = g[30] | (p[30] & g[29]) | (p[30] & p[29] & g[28]) | (p[30] & p[29] & p[28] & g[27]) | (p[30] & p[29] & p[28] & p[27] & g[26]) | (p[30] & p[29] & p[28] & p[27] & p[26] & g[25]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & g[24]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & g[23]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & g[22]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & g[21]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & g[20]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & g[19]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & g[18]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & g[17]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & g[16]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30]);
    assign c[31] = g[31] | (p[31] & g[30]) | (p[31] & p[30] & g[29]) | (p[31] & p[30] & p[29] & g[28]) | (p[31] & p[30] & p[29] & p[28] & g[27]) | (p[31] & p[30] & p[29] & p[28] & p[27] & g[26]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & g[25]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & g[24]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & g[23]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & g[22]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & g[21]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & g[20]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & g[19]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & g[18]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & g[17]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & g[16]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & g[15]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & g[14]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & g[13]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & g[12]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & g[11]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & g[10]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & g[9]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & g[8]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & g[7]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & g[6]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & g[5]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & g[4]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & g[3]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & g[2]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & g[1]) | (p[31] & p[30] & p[29] & p[28] & p[27] & p[26] & p[25] & p[24] & p[23] & p[22] & p[21] & p[20] & p[19] & p[18] & p[17] & p[16] & p[15] & p[14] & p[13] & p[12] & p[11] & p[10] & p[9] & p[8] & p[7] & p[6] & p[5] & p[4] & p[3] & p[2] & p[1] & g[0])| (cin & p[0] & p[1] & p[2] & p[3] & p[4] & p[5] & p[6] & p[7] & p[8] & p[9] & p[10] & p[11] & p[12] & p[13] & p[14] & p[15] & p[16] & p[17] & p[18] & p[19] & p[20] & p[21] & p[22] & p[23] & p[24] & p[25] & p[26] & p[27] & p[28] & p[29] & p[30] & p[31]);
    assign sum[0] = p[0] ^ cin;
    assign sum[1] = p[1] ^ c[0];
    assign sum[2] = p[2] ^ c[1];
    assign sum[3] = p[3] ^ c[2];
    assign sum[4] = p[4] ^ c[3];
    assign sum[5] = p[5] ^ c[4];
    assign sum[6] = p[6] ^ c[5];
    assign sum[7] = p[7] ^ c[6];
    assign sum[8] = p[8] ^ c[7];
    assign sum[9] = p[9] ^ c[8];
    assign sum[10] = p[10] ^ c[9];
    assign sum[11] = p[11] ^ c[10];
    assign sum[12] = p[12] ^ c[11];
    assign sum[13] = p[13] ^ c[12];
    assign sum[14] = p[14] ^ c[13];
    assign sum[15] = p[15] ^ c[14];
    assign sum[16] = p[16] ^ c[15];
    assign sum[17] = p[17] ^ c[16];
    assign sum[18] = p[18] ^ c[17];
    assign sum[19] = p[19] ^ c[18];
    assign sum[20] = p[20] ^ c[19];
    assign sum[21] = p[21] ^ c[20];
    assign sum[22] = p[22] ^ c[21];
    assign sum[23] = p[23] ^ c[22];
    assign sum[24] = p[24] ^ c[23];
    assign sum[25] = p[25] ^ c[24];
    assign sum[26] = p[26] ^ c[25];
    assign sum[27] = p[27] ^ c[26];
    assign sum[28] = p[28] ^ c[27];
    assign sum[29] = p[29] ^ c[28];
    assign sum[30] = p[30] ^ c[29];
    assign sum[31] = p[31] ^ c[30];
    assign Over = c[31];
endmodule

module Shift(input [4:0] shift_bit, input [31:0] B, input[5:0] Op, output [31:0] Result);
    wire [31:0] R_Shift;
    wire [31:0] L_Shift;
    wire [31:0] AR_Shift;
    assign R_Shift = B >> shift_bit;
    assign L_Shift = B << shift_bit;
    assign AR_Shift = $signed(B) >>> shift_bit;
    assign Result =(Op[1])?((Op[0])? AR_Shift : R_Shift):L_Shift;
endmodule

module Logic(input [31:0] A, input [31:0] B, input [5:0] Op, output [31:0] Result);
    wire [31:0] AND_ANS;
    wire [31:0] OR_ANS;
    wire [31:0] XOR_ANS;
    wire [31:0] NOR_ANS;
    assign AND_ANS = A & B;
    assign OR_ANS = A | B;
    assign XOR_ANS = A ^ B;
    assign NOR_ANS = ~(A | B);
    assign Result = (Op[0])?((Op[1])?NOR_ANS:OR_ANS):((Op[1])?XOR_ANS:AND_ANS);
endmodule

module alu(input[31:0] A, input[31:0] B, input[5:0] Op, output[31:0] C, output Over, output zero);
    wire [31:0] mid_B;
    wire [31:0]output_sum;
    wire [31:0]output_shift;
    wire [31:0]output_logic;
    wire [4:0]shift_bit;
    wire [2:0]over; 
    assign shift_bit = A[4:0];
    assign mid_B = (Op[1])? ~B:B;
    Adder_32 Adder_321(A, mid_B, Op[1], output_sum, over[0]);
    Shift Shift1(shift_bit, B, Op, output_shift);
    assign over[1] = 0;
    Logic Logic1(A, B, Op, output_logic);
    assign over[2] = 0;
    assign C = (Op[5])?((Op[2])?output_logic:output_sum):output_shift;
    assign zero = (C[31:0] == 32'b00000000000000000000000000000000)?1:0;
    assign Over = (Op[5])?((Op[2])?over[1]:((~Op[0])&((A[31]==mid_B[31])&(~(A[31]==output_sum[31]))))):over[2]; 
endmodule
